library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity add is
end add;

architecture Behavioral of add is

begin


end Behavioral;

