library ieee;
use ieee.std_logic_1164.all;


entity subtract is
end subtract;

architecture behavioral of subtract is

begin


end behavioral;

