library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity subtract is
end subtract;

architecture Behavioral of subtract is

begin


end Behavioral;

