library ieee;
use ieee.std_logic_1164.all;

entity multiply is
end multiply;

architecture behavioral of multiply is

begin


end behavioral;

