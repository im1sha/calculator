library ieee;
use ieee.std_logic_1164.all;

entity divide is
end divide;

architecture behavioral of divide is

begin


end behavioral;

